// ============================================================================
//   Ver  :| Author					:| Mod. Date :| Changes Made:
//   V1.0 :| viCppDev			   :| 01/02/2021:| Demultiplexor
// ============================================================================

module Demultiplexor (input wire [8:0] dataIN, output wire [8:0] dataOUTA, output wire [8:0] dataOUTB, input wire sel);

	assign dataOUTA = (dataIN)*(!sel);
	assign dataOUTB = (dataIN)*sel;	

endmodule